module app

fn main() {
	println('Hello World!')
}
